----------------------------------------------------------------------------
-- Title : VGA Controller
-- Project : Chip Design BEL4
----------------------------------------------------------------------------
-- File : tb_prescaler_.vhd
-- Author : Resch
-- Company : FHTW
-- Last update: 01.05.2018
-- Platform : VHDL, Modelsim 10.5b, Xilinx Vivado 2016.1
----------------------------------------------------------------------------
-- Description: TESTBENCH ENTITY Prescaler to generate 25MHz signal
----------------------------------------------------------------------------
-- Revisions : 0
-- Date         Version	Author  Description
-- 2018.02.18   0.1     Resch   Projectstart
-- 2018.05.01   0.2     Resch   final code style check and comments
---------------------------------------------------------------------------- 

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity tb_prescaler is

end tb_prescaler;